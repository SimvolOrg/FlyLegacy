<HTML>
<HEAD>
<META HTTP-EQUIV="Content-Type" CONTENT="text/html; charset=windows-1252">
<META NAME="Generator" CONTENT="Microsoft Word 97">
<TITLE>&lt;bgno&gt; ========== BEGIN CAirplane OBJECT ==========</TITLE>
</HEAD>
<BODY>
<FONT FACE="Courier New" SIZE=2><P>&lt;bgno&gt; ========== BEGIN CAirplane OBJECT ==========</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;//</P>
<P>&#9;//&#9;Base Aircraft Info (Fix #1)</P>
<P>&#9;//</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;&lt;mxdt&gt; -- Min Frame Rate (fps)</P>
<P>&#9;35</P>
<P>&#9;&lt;name&gt; -- object name --</P>
<P>&#9;Cessna 172R Skyhawk</P>
<P>&#9;&lt;acid&gt; -- aircraft tail number --</P>
<P>&#9;N234SG</P>
<P>&#9;&lt;make&gt; -- manufacturer (cessna, piper, navajo, hawker, kingair) Used by phrase system</P>
<P>&#9;cessna</P>
<P>&#9;&lt;CLAS&gt; -- classification --</P>
<P>&#9;1</P>
<P>&#9;&lt;USAG&gt; -- usage --</P>
<P>&#9;1</P>
<P>&#9;&lt;emas&gt; -- empty mass --</P>
<P>&#9;49.73</P>
<P>&#9;&lt;maxM&gt; -- max mass --</P>
<P>&#9;76.15</P>
<P>&#9;&lt;mine&gt; ---- momentOfInertia ---- was 1346.0,1967.0,948.0</P>
<P>&#9;350,2000,4000</P>
<P>&#9;&lt;dcen&gt; ---- dynamic center ----</P>
<P>&#9;0,-1.0,1.25</P>
<P>&#9;&lt;iceR&gt; -- Ice Accumulation Rate (hz) --</P>
<P>&#9;0.006</P>
<P>&#9;&lt;CEIL&gt; - ceiling (ft)</P>
<P>&#9;13500</P>
<P>&#9;&lt;043a&gt; - maxCruiseSpeed (kts) -</P>
<P>&#9;123</P>
<P>&#9;&lt;044a&gt; - Approach Speed (kts) -</P>
<P>&#9;80</P>
<P>&#9;&lt;045a&gt; - Best Climb (fpm) -</P>
<P>&#9;500</P>
<P>&#9;&lt;048a&gt; - Never Exceed Speed (kts) - </P>
<P>&#9;163</P>
<P>&#9;&lt;mxCG&gt; - max cg movement (ft) -</P>
<P>&#9;1.0,1.0,-1.0</P>
<P>&#9;&lt;posG&gt; - Positive G Limit (g) -</P>
<P>&#9;3.8</P>
<P>&#9;&lt;negG&gt; - Negative G Limit (g) -</P>
<P>&#9;-1.52</P>
<P>&#9;&lt;stal&gt; -- Simple Stall Speed (ktas) --</P>
<P>&#9;50</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;//</P>
<P>&#9;//&#9;Visual Aircraft Models</P>
<P>&#9;//</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;&lt;mmgr&gt; ---- model manager info ----</P>
<P>&#9;&lt;bgno&gt; ========== BEGIN MODEL MANAGER ==========</P>
<P>&#9;&#9;&lt;mod2&gt; ---- model entry ----</P>
<P>&#9;&#9;comp</P>
<P>&#9;&#9;skyhh.arm</P>
<P>&#9;&#9;200</P>
<P>&#9;&#9;&lt;mod2&gt;</P>
<P>&#9;&#9;comp</P>
<P>&#9;&#9;skyhm.arm</P>
<P>&#9;&#9;60</P>
<P>&#9;&#9;&lt;mod2&gt;</P>
<P>&#9;&#9;comp</P>
<P>&#9;&#9;skyhl.arm</P>
<P>&#9;&#9;20</P>
<P>&#9;&lt;endo&gt; ========== END MODEL MANAGER ==========</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;//</P>
<P>&#9;//&#9;Visual Shadow Models</P>
<P>&#9;//</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;&lt;shdw&gt; ---- shadow info ----</P>
<P>&#9;&lt;bgno&gt; ========== BEGIN OBJECT ==========</P>
<P>&#9;&#9;&lt;modl&gt; ---- shadow model manager ----</P>
<P>&#9;&#9;&lt;bgno&gt; ----</P>
<P>&#9;&#9;&#9;&lt;modl&gt; -- model entry</P>
<P>&#9;&#9;&#9;comp</P>
<P>&#9;&#9;&#9;cessshad.bin</P>
<P>&#9;&#9;&lt;endo&gt; --- </P>
<P>&#9;&lt;endo&gt; ========== END OBJECT ==========</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;//</P>
<P>&#9;//&#9;Cockpit Panels</P>
<P>&#9;//</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;&lt;ckmg&gt; ---- cockpit manager info ----</P>
<P>&#9;&lt;bgno&gt; ========== BEGIN CCOCKPITMANAGER OBJECT ==========</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- forward cockpit entry ----</P>
<P>&#9;&#9;frnt</P>
<P>&#9;&#9;skyhawk0.pnl</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- upper right cockpit entry ----</P>
<P>&#9;&#9;uprt</P>
<P>&#9;&#9;skyhwk10</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- right cockpit entry ----</P>
<P>&#9;&#9;rght</P>
<P>&#9;&#9;skyhwk20</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- lower right cockpit entry ----</P>
<P>&#9;&#9;lwrt</P>
<P>&#9;&#9;skyhwk30</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- backward cockpit entry ----</P>
<P>&#9;&#9;back</P>
<P>&#9;&#9;skyhwk40</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- lower left cockpit entry ----</P>
<P>&#9;&#9;lwlt</P>
<P>&#9;&#9;skyhwk50</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- left cockpit entry ----</P>
<P>&#9;&#9;left</P>
<P>&#9;&#9;skyhwk60</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- upper left cockpit entry ----</P>
<P>&#9;&#9;uplt</P>
<P>&#9;&#9;skyhwk70</P>
<P>&#9;&#9;&lt;ckpt&gt; ---- floor cockpit entry ----</P>
<P>&#9;&#9;floo</P>
<P>&#9;&#9;skyhwk01.pnl</P>
<P>&#9;&lt;endo&gt; ========== END CCOCKPITMANAGER OBJECT ==========</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;//</P>
<P>&#9;//&#9;Mini Cockpit Panel</P>
<P>&#9;//</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;&lt;mini&gt; ---- mini cockpit panel file ----</P>
<P>&#9;miniskyh.pnl</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;//</P>
<P>&#9;//&#9;Available Cameras</P>
<P>&#9;//</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;&lt;cmgr&gt; -- camera manager info --</P>
<P>&#9;&lt;bgno&gt; ========== BEGIN CCAMERAMANAGER OBJECT ==========</P>
<P>&#9;&#9;&lt;came&gt; ---- camera entry ----</P>
<P>&#9;&#9;cock</P>
<P>&#9;&#9;&lt;bgno&gt; ========== BEGIN CCAMERA OBJECT ==========</P>
<P>&#9;&#9;&#9;&lt;seat&gt; ---- seat location (p,b,h,x,y,z) ----</P>
<P>&#9;&#9;&#9;0</P>
<P>&#9;&#9;&#9;0</P>
<P>&#9;&#9;&#9;0</P>
<P>&#9;&#9;&#9;0.0</P>
<P>&#9;&#9;&#9;5.0</P>
<P>&#9;&#9;&#9;4.0</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;frnt</P>
<P>&#9;&#9;&#9;&#9;&lt;main&gt; ---- default ----</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;0.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;uplt</P>
<P>&#9;&#9;&#9;&#9;uprt</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;floo</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;uprt</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;45.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;frnt</P>
<P>&#9;&#9;&#9;&#9;rght</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;rght</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;90.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;uprt</P>
<P>&#9;&#9;&#9;&#9;lwrt</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;lwrt</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;135.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;rght</P>
<P>&#9;&#9;&#9;&#9;back</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;back</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;180.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;lwrt</P>
<P>&#9;&#9;&#9;&#9;lwlt</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;lwlt</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;225.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;back</P>
<P>&#9;&#9;&#9;&#9;left</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;left</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;270.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;lwlt</P>
<P>&#9;&#9;&#9;&#9;uplt</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;uplt</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;315.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;left</P>
<P>&#9;&#9;&#9;&#9;frnt</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&#9;&lt;panl&gt; ---- panel ----</P>
<P>&#9;&#9;&#9;&lt;bgno&gt; ---- begin ----</P>
<P>&#9;&#9;&#9;&#9;&lt;id__&gt; ---- id ----</P>
<P>&#9;&#9;&#9;&#9;floo</P>
<P>&#9;&#9;&#9;&#9;&lt;hdg_&gt; ---- heading ----</P>
<P>&#9;&#9;&#9;&#9;0.0</P>
<P>&#9;&#9;&#9;&#9;&lt;ptch&gt; ---- pitch ----</P>
<P>&#9;&#9;&#9;&#9;45.0</P>
<P>&#9;&#9;&#9;&#9;&lt;pnls&gt; ---- panels (L,R,U,D) ----</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&#9;frnt</P>
<P>&#9;&#9;&#9;&#9;NONE</P>
<P>&#9;&#9;&#9;&lt;endo&gt; ---- end ----</P>
<P>&#9;&#9;&lt;endo&gt; ========== END CCAMERA OBJECT ==========</P>
<P>&#9;&#9;&lt;came&gt; ---- camera entry ----</P>
<P>&#9;&#9;spot</P>
<P>&#9;&#9;&lt;bgno&gt; ========== BEGIN CCAMERA OBJECT ==========</P>
<P>&#9;&#9;&lt;endo&gt; ========== END CCAMERA OBJECT ==========</P>
<P>&#9;&#9;&lt;came&gt; ---- camera entry ----</P>
<P>&#9;&#9;flyb</P>
<P>&#9;&#9;&lt;bgno&gt; ========== BEGIN CCAMERA OBJECT ==========</P>
<P>&#9;&#9;&lt;endo&gt; ========== END CCAMERA OBJECT ==========</P>
<P>&#9;&#9;&lt;came&gt; ---- camera entry ----</P>
<P>&#9;&#9;towr</P>
<P>&#9;&#9;&lt;bgno&gt; ========== BEGIN CCAMERA OBJECT ==========</P>
<P>&#9;&#9;&lt;endo&gt; ========== END CCAMERA OBJECT ==========</P>
<P>&#9;&lt;endo&gt; ========== END CCAMERAMANAGER OBJECT ==========</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;//</P>
<P>&#9;//&#9;Variable Loads</P>
<P>&#9;//</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;&lt;vLdm&gt; - variable Load manager -</P>
<P>&#9;&lt;bgno&gt;</P>
<P>&#9;&#9;&lt;unit&gt; - Single Load Entry -</P>
<P>&#9;&#9;&lt;bgno&gt;</P>
<P>&#9;&#9;&#9;&lt;name&gt; - name of Load -</P>
<P>&#9;&#9;&#9;Pilot</P>
<P>&#9;&#9;&#9;&lt;bPos&gt; - location of load WRT Design CG (fT) -</P>
<P>&#9;&#9;&#9;0,0,0</P>
<P>&#9;&#9;&#9;&lt;load&gt; - weight at load location (lbs) -</P>
<P>&#9;&#9;&#9;170</P>
<P>&#9;&#9;&#9;&lt;hiLm&gt; - max weight limit (lbs) -</P>
<P>&#9;&#9;&#9;300</P>
<P>&#9;&#9;&#9;&lt;uloc&gt; - UI Location</P>
<P>&#9;&#9;&#9;261</P>
<P>&#9;&#9;&#9;290</P>
<P>&#9;&#9;&#9;&lt;utyp&gt; - UI Type Info</P>
<P>&#9;&#9;&#9;Pilot</P>
<P>&#9;&#9;&#9;LW-Pilot.bmp</P>
<P>&#9;&#9;&lt;endo&gt;</P>
<P>&#9;&lt;endo&gt;</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;//</P>
<P>&#9;//&#9;Ground Suspension</P>
<P>&#9;//</P>
<P>&#9;///////////////////////////////////////////////////</P>
<P>&#9;&lt;sspm&gt; ========== Suspension Manager ===========</P>
<P>&#9;&lt;bgno&gt; ========== BEGIN suspension ==========</P>
<P>&#9;&#9;&lt;susp&gt; -- suspension info</P>
<P>&#9;&#9;&lt;bgno&gt; -- begin independent suspension info --</P>
<P>&#9;&#9;&#9;&lt;name&gt; -- wheel part name --</P>
<P>&#9;&#9;&#9;nosewheel</P>
<P>&#9;&#9;&#9;&lt;damn&gt; -- wheel damage region name --</P>
<P>&#9;&#9;&#9;frontSTire</P>
<P>&#9;&#9;&#9;&lt;actn&gt; - strut action -</P>
<P>&#9;&#9;&#9;0</P>
<P>&#9;&#9;&#9;&lt;ster&gt; -- steerable wheel --</P>
<P>&#9;&#9;&#9;1</P>
<P>&#9;&#9;&#9;&lt;mStr&gt; -- max steer angle (deg) --</P>
<P>&#9;&#9;&#9;12.0</P>
<P>&#9;&#9;&#9;&lt;maxC&gt; -- max compression --</P>
<P>&#9;&#9;&#9;0.1</P>
<P>&#9;&#9;&#9;&lt;damR&gt; -- damping ratio --</P>
<P>&#9;&#9;&#9;0.9</P>
<P>&#9;&#9;&lt;endo&gt; -- end independent suspension info --</P>
<P>&#9;&#9;&lt;susp&gt; -- suspension info</P>
<P>&#9;&#9;&lt;bgno&gt; -- begin independent suspension info --</P>
<P>&#9;&#9;&#9;&lt;name&gt; -- wheel part name --</P>
<P>&#9;&#9;&#9;leftwheel</P>
<P>&#9;&#9;&#9;&lt;actn&gt; - beam action -</P>
<P>&#9;&#9;&#9;1</P>
<P>&#9;&#9;&#9;&lt;damn&gt; -- wheel damage region name --</P>
<P>&#9;&#9;&#9;leftBTire</P>
<P>&#9;&#9;&#9;&lt;brak&gt; -- wheel has brake --</P>
<P>&#9;&#9;&#9;-1</P>
<P>&#9;&#9;&#9;&lt;maxC&gt; -- max compression --</P>
<P>&#9;&#9;&#9;0.5</P>
<P>&#9;&#9;&#9;&lt;damR&gt; -- damping ratio --</P>
<P>&#9;&#9;&#9;0.9</P>
<P>&#9;&#9;&lt;endo&gt; -- end independent suspension info --</P>
<P>&#9;&#9;&lt;susp&gt; -- suspension info</P>
<P>&#9;&#9;&lt;bgno&gt; -- begin independent suspension info --</P>
<P>&#9;&#9;&#9;&lt;name&gt; -- wheel part name --</P>
<P>&#9;&#9;&#9;rightwheel</P>
<P>&#9;&#9;&#9;&lt;actn&gt; - beam action -</P>
<P>&#9;&#9;&#9;1</P>
<P>&#9;&#9;&#9;&lt;damn&gt; -- wheel damage region name --</P>
<P>&#9;&#9;&#9;rightBTire</P>
<P>&#9;&#9;&#9;&lt;brak&gt; -- wheel has brake --</P>
<P>&#9;&#9;&#9;1</P>
<P>&#9;&#9;&#9;&lt;maxC&gt; -- max compression --</P>
<P>&#9;&#9;&#9;0.5</P>
<P>&#9;&#9;&#9;&lt;damR&gt; -- damping ratio --</P>
<P>&#9;&#9;&#9;0.9</P>
<P>&#9;&#9;&lt;endo&gt; -- end independent suspension info --</P>
<P>&#9;&lt;endo&gt; ========== END SUSPENSION ==========</P>
<P>&nbsp;</P>
<P>&lt;endo&gt; ========== END CAirplane OBJECT ==========</P>
</FONT></BODY>
</HTML>
